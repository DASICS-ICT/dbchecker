/* =========================================
* Top module wrapper of an accelerator role
*
* Author: Yisong Chang (changyisong@ict.ac.cn)
* Date: 29/01/2021
* Version: v0.0.1
*===========================================
*/

`timescale 10 ns / 1 ns

module dbchecker_wrapper (
  input         clock,
  input         reset,

  input  [31:0] s_axil_ctrl_araddr,
  input  [2:0]  s_axil_ctrl_arprot,
  output        s_axil_ctrl_arready,
  input         s_axil_ctrl_arvalid,
  input  [31:0] s_axil_ctrl_awaddr,
  input  [2:0]  s_axil_ctrl_awprot,
  output        s_axil_ctrl_awready,
  input         s_axil_ctrl_awvalid,
  input         s_axil_ctrl_bready,
  output [1:0]  s_axil_ctrl_bresp,
  output        s_axil_ctrl_bvalid,
  output [31:0] s_axil_ctrl_rdata,
  input         s_axil_ctrl_rready,
  output [1:0]  s_axil_ctrl_rresp,
  output        s_axil_ctrl_rvalid,
  input  [31:0] s_axil_ctrl_wdata,
  output        s_axil_ctrl_wready,
  input  [3:0]  s_axil_ctrl_wstrb,
  input         s_axil_ctrl_wvalid,


  input  [31:0] s_axi_io_tx_araddr,
  input  [1:0]  s_axi_io_tx_arburst,
  input  [3:0]  s_axi_io_tx_arcache,
  input  [7:0]  s_axi_io_tx_arlen,
  input  [0:0]  s_axi_io_tx_arlock,
  input  [2:0]  s_axi_io_tx_arprot,
  input  [3:0]  s_axi_io_tx_arqos,
  input  [3:0]  s_axi_io_tx_arregion,
  output        s_axi_io_tx_arready,
  input  [2:0]  s_axi_io_tx_arsize,
  input         s_axi_io_tx_arvalid,
  input  [31:0] s_axi_io_tx_awaddr,
  input  [1:0]  s_axi_io_tx_awburst,
  input  [3:0]  s_axi_io_tx_awcache,
  input  [7:0]  s_axi_io_tx_awlen,
  input  [0:0]  s_axi_io_tx_awlock,
  input  [2:0]  s_axi_io_tx_awprot,
  input  [3:0]  s_axi_io_tx_awqos,
  input  [3:0]  s_axi_io_tx_awregion,
  output        s_axi_io_tx_awready,
  input  [2:0]  s_axi_io_tx_awsize,
  input         s_axi_io_tx_awvalid,
  input         s_axi_io_tx_bready,
  output [1:0]  s_axi_io_tx_bresp,
  output        s_axi_io_tx_bvalid,
  output [31:0] s_axi_io_tx_rdata,
  output        s_axi_io_tx_rlast,
  input         s_axi_io_tx_rready,
  output [1:0]  s_axi_io_tx_rresp,
  output        s_axi_io_tx_rvalid,
  input  [31:0] s_axi_io_tx_wdata,
  input         s_axi_io_tx_wlast,
  output        s_axi_io_tx_wready,
  input  [15:0] s_axi_io_tx_wstrb,
  input         s_axi_io_tx_wvalid,

  output  [31:0] m_axi_io_tx_araddr,
  output  [1:0]  m_axi_io_tx_arburst,
  output  [3:0]  m_axi_io_tx_arcache,
  output  [7:0]  m_axi_io_tx_arlen,
  output  [0:0]  m_axi_io_tx_arlock,
  output  [2:0]  m_axi_io_tx_arprot,
  output  [3:0]  m_axi_io_tx_arqos,
  input          m_axi_io_tx_arready,
  output  [2:0]  m_axi_io_tx_arsize,
  output         m_axi_io_tx_arvalid,
  output  [31:0] m_axi_io_tx_awaddr,
  output  [1:0]  m_axi_io_tx_awburst,
  output  [3:0]  m_axi_io_tx_awcache,
  output  [7:0]  m_axi_io_tx_awlen,
  output  [0:0]  m_axi_io_tx_awlock,
  output  [2:0]  m_axi_io_tx_awprot,
  output  [3:0]  m_axi_io_tx_awqos,
  input          m_axi_io_tx_awready,
  output  [2:0]  m_axi_io_tx_awsize,
  output         m_axi_io_tx_awvalid,
  output         m_axi_io_tx_bready,
  input   [1:0]  m_axi_io_tx_bresp,
  input          m_axi_io_tx_bvalid,
  input   [31:0] m_axi_io_tx_rdata,
  input          m_axi_io_tx_rlast,
  output         m_axi_io_tx_rready,
  input   [1:0]  m_axi_io_tx_rresp,
  input          m_axi_io_tx_rvalid,
  output  [31:0] m_axi_io_tx_wdata,
  output         m_axi_io_tx_wlast,
  input          m_axi_io_tx_wready,
  output  [15:0] m_axi_io_tx_wstrb,
  output         m_axi_io_tx_wvalid,

  input  [63:0] s_axi_io_rx_araddr,
  input  [1:0]  s_axi_io_rx_arburst,
  input  [3:0]  s_axi_io_rx_arcache,
  input  [7:0]  s_axi_io_rx_arlen,
  input  [0:0]  s_axi_io_rx_arlock,
  input  [2:0]  s_axi_io_rx_arprot,
  input  [3:0]  s_axi_io_rx_arqos,
  input  [3:0]  s_axi_io_rx_arregion,
  output        s_axi_io_rx_arready,
  input  [2:0]  s_axi_io_rx_arsize,
  input         s_axi_io_rx_arvalid,
  input  [63:0] s_axi_io_rx_awaddr,
  input  [1:0]  s_axi_io_rx_awburst,
  input  [3:0]  s_axi_io_rx_awcache,
  input  [7:0]  s_axi_io_rx_awlen,
  input  [0:0]  s_axi_io_rx_awlock,
  input  [2:0]  s_axi_io_rx_awprot,
  input  [3:0]  s_axi_io_rx_awqos,
  input  [3:0]  s_axi_io_rx_awregion,
  output        s_axi_io_rx_awready,
  input  [2:0]  s_axi_io_rx_awsize,
  input         s_axi_io_rx_awvalid,
  input         s_axi_io_rx_bready,
  output [1:0]  s_axi_io_rx_bresp,
  output        s_axi_io_rx_bvalid,
  output [127:0]s_axi_io_rx_rdata,
  output        s_axi_io_rx_rlast,
  input         s_axi_io_rx_rready,
  output [1:0]  s_axi_io_rx_rresp,
  output        s_axi_io_rx_rvalid,
  input  [127:0]s_axi_io_rx_wdata,
  input         s_axi_io_rx_wlast,
  output        s_axi_io_rx_wready,
  input  [15:0] s_axi_io_rx_wstrb,
  input         s_axi_io_rx_wvalid,

  output  [35:0] m_axi_io_rx_araddr,
  output  [1:0]  m_axi_io_rx_arburst,
  output  [3:0]  m_axi_io_rx_arcache,
  output  [7:0]  m_axi_io_rx_arlen,
  output  [0:0]  m_axi_io_rx_arlock,
  output  [2:0]  m_axi_io_rx_arprot,
  output  [3:0]  m_axi_io_rx_arqos,
  input          m_axi_io_rx_arready,
  output  [2:0]  m_axi_io_rx_arsize,
  output         m_axi_io_rx_arvalid,
  output  [35:0] m_axi_io_rx_awaddr,
  output  [1:0]  m_axi_io_rx_awburst,
  output  [3:0]  m_axi_io_rx_awcache,
  output  [7:0]  m_axi_io_rx_awlen,
  output  [0:0]  m_axi_io_rx_awlock,
  output  [2:0]  m_axi_io_rx_awprot,
  output  [3:0]  m_axi_io_rx_awqos,
  input          m_axi_io_rx_awready,
  output  [2:0]  m_axi_io_rx_awsize,
  output         m_axi_io_rx_awvalid,
  output         m_axi_io_rx_bready,
  input   [1:0]  m_axi_io_rx_bresp,
  input          m_axi_io_rx_bvalid,
  input   [127:0]m_axi_io_rx_rdata,
  input          m_axi_io_rx_rlast,
  output         m_axi_io_rx_rready,
  input   [1:0]  m_axi_io_rx_rresp,
  input          m_axi_io_rx_rvalid,
  output  [127:0]m_axi_io_rx_wdata,
  output         m_axi_io_rx_wlast,
  input          m_axi_io_rx_wready,
  output  [15:0] m_axi_io_rx_wstrb,
  output         m_axi_io_rx_wvalid

);

DBChecker DBChecker_0(
  .clock(clock),
  .reset(reset),

  .s_axil_ctrl_ar_bits_addr(s_axil_ctrl_araddr),
  .s_axil_ctrl_ar_bits_prot(s_axil_ctrl_arprot),
  .s_axil_ctrl_ar_ready(s_axil_ctrl_arready),
  .s_axil_ctrl_ar_valid(s_axil_ctrl_arvalid),
  .s_axil_ctrl_aw_bits_addr(s_axil_ctrl_awaddr),
  .s_axil_ctrl_aw_bits_prot(s_axil_ctrl_awprot),
  .s_axil_ctrl_aw_ready(s_axil_ctrl_awready),
  .s_axil_ctrl_aw_valid(s_axil_ctrl_awvalid),
  .s_axil_ctrl_b_ready(s_axil_ctrl_bready),
  .s_axil_ctrl_b_bits_resp(s_axil_ctrl_bresp),
  .s_axil_ctrl_b_valid(s_axil_ctrl_bvalid),
  .s_axil_ctrl_r_bits_data(s_axil_ctrl_rdata),
  .s_axil_ctrl_r_ready(s_axil_ctrl_rready),
  .s_axil_ctrl_r_bits_resp(s_axil_ctrl_rresp),
  .s_axil_ctrl_r_valid(s_axil_ctrl_rvalid),
  .s_axil_ctrl_w_bits_data(s_axil_ctrl_wdata),
  .s_axil_ctrl_w_ready(s_axil_ctrl_wready),
  .s_axil_ctrl_w_bits_strb(s_axil_ctrl_wstrb),
  .s_axil_ctrl_w_valid(s_axil_ctrl_wvalid),
  
  .s_axi_io_tx_ar_bits_addr(s_axi_io_tx_araddr),
  .s_axi_io_tx_ar_bits_burst(s_axi_io_tx_arburst),
  .s_axi_io_tx_ar_bits_cache(s_axi_io_tx_arcache),
  .s_axi_io_tx_ar_bits_len(s_axi_io_tx_arlen),
  .s_axi_io_tx_ar_bits_lock(s_axi_io_tx_arlock),
  .s_axi_io_tx_ar_bits_prot(s_axi_io_tx_arprot),
  .s_axi_io_tx_ar_bits_qos(s_axi_io_tx_arqos),
  .s_axi_io_tx_ar_ready(s_axi_io_tx_arready),
  .s_axi_io_tx_ar_bits_size(s_axi_io_tx_arsize),
  .s_axi_io_tx_ar_valid(s_axi_io_tx_arvalid),
  .s_axi_io_tx_aw_bits_addr(s_axi_io_tx_awaddr),
  .s_axi_io_tx_aw_bits_burst(s_axi_io_tx_awburst),
  .s_axi_io_tx_aw_bits_cache(s_axi_io_tx_awcache),
  .s_axi_io_tx_aw_bits_len(s_axi_io_tx_awlen),
  .s_axi_io_tx_aw_bits_lock(s_axi_io_tx_awlock),
  .s_axi_io_tx_aw_bits_prot(s_axi_io_tx_awprot),
  .s_axi_io_tx_aw_bits_qos(s_axi_io_tx_awqos),
  .s_axi_io_tx_aw_ready(s_axi_io_tx_awready),
  .s_axi_io_tx_aw_bits_size(s_axi_io_tx_awsize),
  .s_axi_io_tx_aw_valid(s_axi_io_tx_awvalid),
  .s_axi_io_tx_b_ready(s_axi_io_tx_bready),
  .s_axi_io_tx_b_bits_resp(s_axi_io_tx_bresp),
  .s_axi_io_tx_b_valid(s_axi_io_tx_bvalid),
  .s_axi_io_tx_r_bits_data(s_axi_io_tx_rdata),
  .s_axi_io_tx_r_bits_last(s_axi_io_tx_rlast),
  .s_axi_io_tx_r_ready(s_axi_io_tx_rready),
  .s_axi_io_tx_r_bits_resp(s_axi_io_tx_rresp),
  .s_axi_io_tx_r_valid(s_axi_io_tx_rvalid),
  .s_axi_io_tx_w_bits_data(s_axi_io_tx_wdata),
  .s_axi_io_tx_w_bits_last(s_axi_io_tx_wlast),
  .s_axi_io_tx_w_ready(s_axi_io_tx_wready),
  .s_axi_io_tx_w_bits_strb(s_axi_io_tx_wstrb),
  .s_axi_io_tx_w_valid(s_axi_io_tx_wvalid),

  .m_axi_io_tx_ar_bits_addr(m_axi_io_tx_araddr),
  .m_axi_io_tx_ar_bits_burst(m_axi_io_tx_arburst),
  .m_axi_io_tx_ar_bits_cache(m_axi_io_tx_arcache),
  .m_axi_io_tx_ar_bits_len(m_axi_io_tx_arlen),
  .m_axi_io_tx_ar_bits_lock(m_axi_io_tx_arlock),
  .m_axi_io_tx_ar_bits_prot(m_axi_io_tx_arprot),
  .m_axi_io_tx_ar_bits_qos(m_axi_io_tx_arqos),
  .m_axi_io_tx_ar_bits_region(m_axi_io_tx_arregion),
  .m_axi_io_tx_ar_ready(m_axi_io_tx_arready),
  .m_axi_io_tx_ar_bits_size(m_axi_io_tx_arsize),
  .m_axi_io_tx_ar_valid(m_axi_io_tx_arvalid),
  .m_axi_io_tx_aw_bits_addr(m_axi_io_tx_awaddr),
  .m_axi_io_tx_aw_bits_burst(m_axi_io_tx_awburst),
  .m_axi_io_tx_aw_bits_cache(m_axi_io_tx_awcache),
  .m_axi_io_tx_aw_bits_len(m_axi_io_tx_awlen),
  .m_axi_io_tx_aw_bits_lock(m_axi_io_tx_awlock),
  .m_axi_io_tx_aw_bits_prot(m_axi_io_tx_awprot),
  .m_axi_io_tx_aw_bits_qos(m_axi_io_tx_awqos),
  .m_axi_io_tx_aw_bits_region(m_axi_io_tx_awregion),
  .m_axi_io_tx_aw_ready(m_axi_io_tx_awready),
  .m_axi_io_tx_aw_bits_size(m_axi_io_tx_awsize),
  .m_axi_io_tx_aw_valid(m_axi_io_tx_awvalid),
  .m_axi_io_tx_b_ready(m_axi_io_tx_bready),
  .m_axi_io_tx_b_bits_resp(m_axi_io_tx_bresp),
  .m_axi_io_tx_b_valid(m_axi_io_tx_bvalid),
  .m_axi_io_tx_r_bits_data(m_axi_io_tx_rdata),
  .m_axi_io_tx_r_bits_last(m_axi_io_tx_rlast),
  .m_axi_io_tx_r_ready(m_axi_io_tx_rready),
  .m_axi_io_tx_r_bits_resp(m_axi_io_tx_rresp),
  .m_axi_io_tx_r_valid(m_axi_io_tx_rvalid),
  .m_axi_io_tx_w_bits_data(m_axi_io_tx_wdata),
  .m_axi_io_tx_w_bits_last(m_axi_io_tx_wlast),
  .m_axi_io_tx_w_ready(m_axi_io_tx_wready),
  .m_axi_io_tx_w_bits_strb(m_axi_io_tx_wstrb),
  .m_axi_io_tx_w_valid(m_axi_io_tx_wvalid),

    .s_axi_io_rx_ar_bits_addr(s_axi_io_rx_araddr),
  .s_axi_io_rx_ar_bits_burst(s_axi_io_rx_arburst),
  .s_axi_io_rx_ar_bits_cache(s_axi_io_rx_arcache),
  .s_axi_io_rx_ar_bits_len(s_axi_io_rx_arlen),
  .s_axi_io_rx_ar_bits_lock(s_axi_io_rx_arlock),
  .s_axi_io_rx_ar_bits_prot(s_axi_io_rx_arprot),
  .s_axi_io_rx_ar_bits_qos(s_axi_io_rx_arqos),
  .s_axi_io_rx_ar_ready(s_axi_io_rx_arready),
  .s_axi_io_rx_ar_bits_size(s_axi_io_rx_arsize),
  .s_axi_io_rx_ar_valid(s_axi_io_rx_arvalid),
  .s_axi_io_rx_aw_bits_addr(s_axi_io_rx_awaddr),
  .s_axi_io_rx_aw_bits_burst(s_axi_io_rx_awburst),
  .s_axi_io_rx_aw_bits_cache(s_axi_io_rx_awcache),
  .s_axi_io_rx_aw_bits_len(s_axi_io_rx_awlen),
  .s_axi_io_rx_aw_bits_lock(s_axi_io_rx_awlock),
  .s_axi_io_rx_aw_bits_prot(s_axi_io_rx_awprot),
  .s_axi_io_rx_aw_bits_qos(s_axi_io_rx_awqos),
  .s_axi_io_rx_aw_ready(s_axi_io_rx_awready),
  .s_axi_io_rx_aw_bits_size(s_axi_io_rx_awsize),
  .s_axi_io_rx_aw_valid(s_axi_io_rx_awvalid),
  .s_axi_io_rx_b_ready(s_axi_io_rx_bready),
  .s_axi_io_rx_b_bits_resp(s_axi_io_rx_bresp),
  .s_axi_io_rx_b_valid(s_axi_io_rx_bvalid),
  .s_axi_io_rx_r_bits_data(s_axi_io_rx_rdata),
  .s_axi_io_rx_r_bits_last(s_axi_io_rx_rlast),
  .s_axi_io_rx_r_ready(s_axi_io_rx_rready),
  .s_axi_io_rx_r_bits_resp(s_axi_io_rx_rresp),
  .s_axi_io_rx_r_valid(s_axi_io_rx_rvalid),
  .s_axi_io_rx_w_bits_data(s_axi_io_rx_wdata),
  .s_axi_io_rx_w_bits_last(s_axi_io_rx_wlast),
  .s_axi_io_rx_w_ready(s_axi_io_rx_wready),
  .s_axi_io_rx_w_bits_strb(s_axi_io_rx_wstrb),
  .s_axi_io_rx_w_valid(s_axi_io_rx_wvalid),

  .m_axi_io_rx_ar_bits_addr(m_axi_io_rx_araddr),
  .m_axi_io_rx_ar_bits_burst(m_axi_io_rx_arburst),
  .m_axi_io_rx_ar_bits_cache(m_axi_io_rx_arcache),
  .m_axi_io_rx_ar_bits_len(m_axi_io_rx_arlen),
  .m_axi_io_rx_ar_bits_lock(m_axi_io_rx_arlock),
  .m_axi_io_rx_ar_bits_prot(m_axi_io_rx_arprot),
  .m_axi_io_rx_ar_bits_qos(m_axi_io_rx_arqos),
  .m_axi_io_rx_ar_bits_region(m_axi_io_rx_arregion),
  .m_axi_io_rx_ar_ready(m_axi_io_rx_arready),
  .m_axi_io_rx_ar_bits_size(m_axi_io_rx_arsize),
  .m_axi_io_rx_ar_valid(m_axi_io_rx_arvalid),
  .m_axi_io_rx_aw_bits_addr(m_axi_io_rx_awaddr),
  .m_axi_io_rx_aw_bits_burst(m_axi_io_rx_awburst),
  .m_axi_io_rx_aw_bits_cache(m_axi_io_rx_awcache),
  .m_axi_io_rx_aw_bits_len(m_axi_io_rx_awlen),
  .m_axi_io_rx_aw_bits_lock(m_axi_io_rx_awlock),
  .m_axi_io_rx_aw_bits_prot(m_axi_io_rx_awprot),
  .m_axi_io_rx_aw_bits_qos(m_axi_io_rx_awqos),
  .m_axi_io_rx_aw_bits_region(m_axi_io_rx_awregion),
  .m_axi_io_rx_aw_ready(m_axi_io_rx_awready),
  .m_axi_io_rx_aw_bits_size(m_axi_io_rx_awsize),
  .m_axi_io_rx_aw_valid(m_axi_io_rx_awvalid),
  .m_axi_io_rx_b_ready(m_axi_io_rx_bready),
  .m_axi_io_rx_b_bits_resp(m_axi_io_rx_bresp),
  .m_axi_io_rx_b_valid(m_axi_io_rx_bvalid),
  .m_axi_io_rx_r_bits_data(m_axi_io_rx_rdata),
  .m_axi_io_rx_r_bits_last(m_axi_io_rx_rlast),
  .m_axi_io_rx_r_ready(m_axi_io_rx_rready),
  .m_axi_io_rx_r_bits_resp(m_axi_io_rx_rresp),
  .m_axi_io_rx_r_valid(m_axi_io_rx_rvalid),
  .m_axi_io_rx_w_bits_data(m_axi_io_rx_wdata),
  .m_axi_io_rx_w_bits_last(m_axi_io_rx_wlast),
  .m_axi_io_rx_w_ready(m_axi_io_rx_wready),
  .m_axi_io_rx_w_bits_strb(m_axi_io_rx_wstrb),
  .m_axi_io_rx_w_valid(m_axi_io_rx_wvalid)

);

endmodule
